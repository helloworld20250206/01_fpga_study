library verilog;
use verilog.vl_types.all;
entity top_fpga_vlg_tst is
end top_fpga_vlg_tst;
